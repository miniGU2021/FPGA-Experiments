library verilog;
use verilog.vl_types.all;
entity stb2_59_vlg_sample_tst is
    port(
        CLK_59          : in     vl_logic;
        R_59            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end stb2_59_vlg_sample_tst;
