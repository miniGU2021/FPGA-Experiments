library verilog;
use verilog.vl_types.all;
entity stb2_59_vlg_check_tst is
    port(
        P_59            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end stb2_59_vlg_check_tst;
