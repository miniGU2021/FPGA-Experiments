library verilog;
use verilog.vl_types.all;
entity segsel_59_vlg_vec_tst is
end segsel_59_vlg_vec_tst;
