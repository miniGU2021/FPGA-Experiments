library verilog;
use verilog.vl_types.all;
entity cnt_m10_vlg_vec_tst is
end cnt_m10_vlg_vec_tst;
