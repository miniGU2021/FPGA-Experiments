library verilog;
use verilog.vl_types.all;
entity dynamic_display_m100_vlg_vec_tst is
end dynamic_display_m100_vlg_vec_tst;
