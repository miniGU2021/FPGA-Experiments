library verilog;
use verilog.vl_types.all;
entity stb2_59_vlg_vec_tst is
end stb2_59_vlg_vec_tst;
