library verilog;
use verilog.vl_types.all;
entity cnt6_vlg_sample_tst is
    port(
        p_59            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt6_vlg_sample_tst;
