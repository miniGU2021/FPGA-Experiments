library verilog;
use verilog.vl_types.all;
entity display_vlg_check_tst is
    port(
        DIGOUT_59       : in     vl_logic_vector(7 downto 0);
        SEGOUT_59       : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end display_vlg_check_tst;
