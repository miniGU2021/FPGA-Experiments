library verilog;
use verilog.vl_types.all;
entity cnt_m10_vlg_sample_tst is
    port(
        CLK_59          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt_m10_vlg_sample_tst;
