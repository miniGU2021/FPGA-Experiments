library verilog;
use verilog.vl_types.all;
entity fre_div_59_vlg_sample_tst is
    port(
        CI              : in     vl_logic;
        TI              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end fre_div_59_vlg_sample_tst;
