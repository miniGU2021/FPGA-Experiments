library verilog;
use verilog.vl_types.all;
entity m100_59 is
    port(
        CO              : out    vl_logic;
        CI              : in     vl_logic
    );
end m100_59;
