library verilog;
use verilog.vl_types.all;
entity m100_59_vlg_check_tst is
    port(
        CO              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end m100_59_vlg_check_tst;
