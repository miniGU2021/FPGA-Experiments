library verilog;
use verilog.vl_types.all;
entity digsel_59_vlg_check_tst is
    port(
        DIGOUT_59       : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end digsel_59_vlg_check_tst;
