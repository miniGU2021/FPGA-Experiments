library verilog;
use verilog.vl_types.all;
entity fre_div_59 is
    port(
        CO1             : out    vl_logic;
        CI              : in     vl_logic;
        CO2             : out    vl_logic;
        CO3             : out    vl_logic
    );
end fre_div_59;
