library verilog;
use verilog.vl_types.all;
entity segsel_59_vlg_check_tst is
    port(
        SEGOUT_59       : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end segsel_59_vlg_check_tst;
