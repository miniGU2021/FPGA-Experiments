library verilog;
use verilog.vl_types.all;
entity digsel_vlg_vec_tst is
end digsel_vlg_vec_tst;
