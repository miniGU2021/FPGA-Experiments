library verilog;
use verilog.vl_types.all;
entity cnt6 is
    port(
        Q               : out    vl_logic;
        p_59            : in     vl_logic;
        q_59            : out    vl_logic_vector(3 downto 0)
    );
end cnt6;
