library verilog;
use verilog.vl_types.all;
entity decoder_59_vlg_check_tst is
    port(
        S_59            : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end decoder_59_vlg_check_tst;
