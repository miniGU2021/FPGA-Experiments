library verilog;
use verilog.vl_types.all;
entity cnt_m10 is
    port(
        D_59            : out    vl_logic_vector(3 downto 0);
        CLK_59          : in     vl_logic
    );
end cnt_m10;
