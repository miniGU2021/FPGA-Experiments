library verilog;
use verilog.vl_types.all;
entity stb2_59 is
    port(
        P_59            : out    vl_logic;
        CLK_59          : in     vl_logic;
        R_59            : in     vl_logic
    );
end stb2_59;
