library verilog;
use verilog.vl_types.all;
entity decoder_59 is
    port(
        S_59            : out    vl_logic_vector(6 downto 0);
        D_59            : in     vl_logic_vector(3 downto 0)
    );
end decoder_59;
