library verilog;
use verilog.vl_types.all;
entity fre_div_59_vlg_check_tst is
    port(
        CO1             : in     vl_logic;
        CO2             : in     vl_logic;
        CO3             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fre_div_59_vlg_check_tst;
