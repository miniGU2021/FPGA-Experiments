library verilog;
use verilog.vl_types.all;
entity digsel_59_vlg_vec_tst is
end digsel_59_vlg_vec_tst;
