library verilog;
use verilog.vl_types.all;
entity m100_59_vlg_vec_tst is
end m100_59_vlg_vec_tst;
