library verilog;
use verilog.vl_types.all;
entity decoder_59_vlg_vec_tst is
end decoder_59_vlg_vec_tst;
